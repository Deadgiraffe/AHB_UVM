package pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "seqItem.sv"
    `include "sequence.sv"
    `include "seqr.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "scoreboard.sv"
    `include "env.sv"
    `include "test.sv"

endpackage